***** Spice Netlist for Cell 'Lab9_inv' *****

************** Module Lab9_inv **************
.subckt Lab9_inv vin vout
m1 vout vin gnd gnd scmosn w='0.6u' l='0.4u' m='1' 
m2 vout vin vdd vdd scmosp w='0.6u' l='0.4u' m='1' 
.ends Lab9_inv


.end

