magic
tech scmos
timestamp 1623065174
<< nwell >>
rect -21 0 22 27
<< ntransistor >>
rect -1 -12 1 -7
<< ptransistor >>
rect -1 6 1 16
<< ndiffusion >>
rect -6 -12 -1 -7
rect 1 -12 7 -7
<< pdiffusion >>
rect -6 6 -1 16
rect 1 6 7 16
<< ndcontact >>
rect -10 -12 -6 -7
rect 7 -12 11 -7
<< pdcontact >>
rect -10 6 -6 16
rect 7 6 11 16
<< psubstratepcontact >>
rect -10 -21 -6 -16
rect 7 -21 11 -16
<< nsubstratencontact >>
rect -10 20 -6 24
rect 7 20 11 24
<< polysilicon >>
rect -1 16 1 18
rect -1 -7 1 6
rect -1 -14 1 -12
<< polycontact >>
rect -5 -3 -1 1
<< metal1 >>
rect -6 20 7 24
rect -10 19 11 20
rect -10 16 -6 19
rect -7 -3 -5 1
rect -1 -3 1 0
rect 7 -7 11 6
rect -10 -15 -6 -12
rect -10 -16 11 -15
rect -6 -21 7 -16
<< labels >>
rlabel metal1 -10 -15 -10 -15 1 Gnd
rlabel metal1 8 0 8 0 1 out
rlabel metal1 -9 20 -9 20 5 Vdd
rlabel polycontact -3 -2 -3 -2 1 in
<< end >>
